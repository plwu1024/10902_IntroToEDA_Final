module top (a, b, c, o1);
input a, b, c;
output o1;
wire a, b, c, o1;
and g1 (o1, a, b, c);
endmodule