module top(o, a);
output o;
input a, b, c;
wire t_0, o1; 
and g1(o1, a, b, c);
assign o = t_0;
endmodule
