module top(o, a, b, c);
input a, b, c;
output o;
wire n1;
and g1(o, a, b, c);
endmodule